
module embedded_system (
	clk_clk,
	resetn_reset_n,
	to_hex_readdata);	

	input		clk_clk;
	input		resetn_reset_n;
	output	[31:0]	to_hex_readdata;
endmodule
